// A simple demo of animation, VGA signal generation, and a rotation effect.
// Brandon Pelfrey
// Video at https://www.youtube.com/watch?v=Q7v7Moh8ltM
//
// I'm new to verilog. This code is probably awful.

module top(
  input clk25,   // Onboard 12Mhz Oscillator
  output r0,      // 1-bit VGA Red/Green/Blue
  output g0,
  output b0,
  output hsync,   // VGA H-Sync Signal
  output vsync);  // VGA V-Sync Signal

// VGA has a pixel clock which defines the time between 
// each consecutive pixel. For a given video mode, which is
// 640 x 480 @ 60 fps here, you need a specific pixel clock
// speed. In this case, 25.175 MHz. 'icepll -o 25.175' will
// determine the best coefficients in the PLL equation to
// get as close to this as possible (monitor is pretty
// tolerant to be slightly off).
/*
SB_PLL40_PAD #(
  .FEEDBACK_PATH("SIMPLE"),
  .DIVR(4'b0000),
  .DIVF(7'b1000010),
  .DIVQ(3'b101),
  .FILTER_RANGE(3'b001)
) uut (
  .RESETB(1'b1),
  .BYPASS(1'b0),
  .PACKAGEPIN(clk_in),
  .PLLOUTCORE(clk_out)

);
*/

// Some other constants for the VGA signal. Each line begins
// with actual image data, then an H-Sync front porch, pulse,
// and back porch, which are used for locking onto a signal at
// the monitor. A similar thing happens after the last line
// of color data: There are several lines forming a V-Sync
// front porch, pulse, and back porch.
parameter res_x = 640;
parameter res_y = 480;

parameter hfp = 16;      // horizontal front porch
parameter hpulse = 96;   // hsync pulse length
parameter hbp = 48;      // horizontal back porch

parameter vfp = 10;      // vertical front porch
parameter vpulse = 2;    // vsync pulse length
parameter vbp = 33;      // vertical back porch

parameter hpixels = res_x + hfp + hpulse + hbp; // horizontal pixels per line
parameter vlines  = res_y + vfp + vpulse + vbp; // vertical lines per frame

// Tiled image bitmap which composes the background image.
reg[0:7] tile_data[0:7];

// Some sine wave data which is indexed by position and frame number to
// produce distortions in how the tile data is indexed. The effect is that
// the tile data appears to move on screen, when in fact, the indexing is
// just being manipulated.
reg[7:0] line_shifts[63:0];

initial begin
  tile_data[0] <= 8'b10000001;
  tile_data[1] <= 8'b01000010;
  tile_data[2] <= 8'b00100100;
  tile_data[3] <= 8'b00011100;
  tile_data[4] <= 8'b00011000;
  tile_data[5] <= 8'b00100100;
  tile_data[6] <= 8'b01000010;
  tile_data[7] <= 8'b10000001;

  line_shifts[0] <= 8'd8;
  line_shifts[1] <= 8'd8;
  line_shifts[2] <= 8'd9;
  line_shifts[3] <= 8'd10;
  line_shifts[4] <= 8'd11;
  line_shifts[5] <= 8'd11;
  line_shifts[6] <= 8'd12;
  line_shifts[7] <= 8'd13;
  line_shifts[8] <= 8'd13;
  line_shifts[9] <= 8'd14;
  line_shifts[10] <= 8'd14;
  line_shifts[11] <= 8'd15;
  line_shifts[12] <= 8'd15;
  line_shifts[13] <= 8'd15;
  line_shifts[14] <= 8'd15;
  line_shifts[15] <= 8'd15;
  line_shifts[16] <= 8'd15;
  line_shifts[17] <= 8'd15;
  line_shifts[18] <= 8'd15;
  line_shifts[19] <= 8'd15;
  line_shifts[20] <= 8'd15;
  line_shifts[21] <= 8'd14;
  line_shifts[22] <= 8'd14;
  line_shifts[23] <= 8'd13;
  line_shifts[24] <= 8'd13;
  line_shifts[25] <= 8'd12;
  line_shifts[26] <= 8'd12;
  line_shifts[27] <= 8'd11;
  line_shifts[28] <= 8'd10;
  line_shifts[29] <= 8'd9;
  line_shifts[30] <= 8'd9;
  line_shifts[31] <= 8'd8;
  line_shifts[32] <= 8'd7;
  line_shifts[33] <= 8'd6;
  line_shifts[34] <= 8'd6;
  line_shifts[35] <= 8'd5;
  line_shifts[36] <= 8'd4;
  line_shifts[37] <= 8'd3;
  line_shifts[38] <= 8'd3;
  line_shifts[39] <= 8'd2;
  line_shifts[40] <= 8'd2;
  line_shifts[41] <= 8'd1;
  line_shifts[42] <= 8'd1;
  line_shifts[43] <= 8'd0;
  line_shifts[44] <= 8'd0;
  line_shifts[45] <= 8'd0;
  line_shifts[46] <= 8'd0;
  line_shifts[47] <= 8'd0;
  line_shifts[48] <= 8'd0;
  line_shifts[49] <= 8'd0;
  line_shifts[50] <= 8'd0;
  line_shifts[51] <= 8'd0;
  line_shifts[52] <= 8'd0;
  line_shifts[53] <= 8'd1;
  line_shifts[54] <= 8'd1;
  line_shifts[55] <= 8'd2;
  line_shifts[56] <= 8'd2;
  line_shifts[57] <= 8'd3;
  line_shifts[58] <= 8'd4;
  line_shifts[59] <= 8'd4;
  line_shifts[60] <= 8'd5;
  line_shifts[61] <= 8'd6;
  line_shifts[62] <= 8'd7;
  line_shifts[63] <= 8'd7;
end

// These are our horizontal and vertical positions on
// the screen at any moment (including fp/pulse/bp)
reg [12:0] pix_x;
reg [12:0] pix_y;

// Some state used to compute shifting for the tile data.
reg pix_reg;
reg[8:0] shift_x;
reg[5:0] shift_x_index;
reg[8:0] shift_y;
reg[5:0] shift_y_index;

// Which frame we're on. Used in animation.
reg[15:0] frame_counter = 0;

///////////////////////////////////////////////////////

// The image is rotated by computing rotated positions
//
// --- x' = c*x - s*y
// --- y' = s*x + c*y
//
// where c = cos(theta), s = sin(theta), and theta changes
// each frame.
//
// To avoid multiplication, these equations are mutliplied
// by B=2^k.
//
// --- B*x' = (B*c)*x - (B*s)*y
// --- B*y' = (B*s)*x + (B*c)*y
//
// We can avoid the multiply by simply keeping a running
// sum of each of B*c*x, B*s*y, B*s*x, and B*c*y. This way
// we only need to add constants as we advance the pixel
// one pixel to the right or one line down.
//
// When you need to know the actual (x',y'), you simply
// divide by B, but that's just a power of 2, so do an
// arithmetic right shift by k.
//

// cos(theta) and sin(theta) for 1024 divisions of a single
// rotation. Computed in a little python script.
reg signed[12:0] Cp[1023:0];
reg signed[12:0] Sp[1023:0];

initial begin
Cp[0] <= 11'd1024; Sp[0] <= 11'd0;
Cp[1] <= 11'd1023; Sp[1] <= 11'd6;
Cp[2] <= 11'd1023; Sp[2] <= 11'd12;
Cp[3] <= 11'd1023; Sp[3] <= 11'd18;
Cp[4] <= 11'd1023; Sp[4] <= 11'd25;
Cp[5] <= 11'd1023; Sp[5] <= 11'd31;
Cp[6] <= 11'd1023; Sp[6] <= 11'd37;
Cp[7] <= 11'd1023; Sp[7] <= 11'd44;
Cp[8] <= 11'd1022; Sp[8] <= 11'd50;
Cp[9] <= 11'd1022; Sp[9] <= 11'd56;
Cp[10] <= 11'd1022; Sp[10] <= 11'd62;
Cp[11] <= 11'd1021; Sp[11] <= 11'd69;
Cp[12] <= 11'd1021; Sp[12] <= 11'd75;
Cp[13] <= 11'd1020; Sp[13] <= 11'd81;
Cp[14] <= 11'd1020; Sp[14] <= 11'd87;
Cp[15] <= 11'd1019; Sp[15] <= 11'd94;
Cp[16] <= 11'd1019; Sp[16] <= 11'd100;
Cp[17] <= 11'd1018; Sp[17] <= 11'd106;
Cp[18] <= 11'd1017; Sp[18] <= 11'd112;
Cp[19] <= 11'd1017; Sp[19] <= 11'd119;
Cp[20] <= 11'd1016; Sp[20] <= 11'd125;
Cp[21] <= 11'd1015; Sp[21] <= 11'd131;
Cp[22] <= 11'd1014; Sp[22] <= 11'd137;
Cp[23] <= 11'd1013; Sp[23] <= 11'd144;
Cp[24] <= 11'd1012; Sp[24] <= 11'd150;
Cp[25] <= 11'd1011; Sp[25] <= 11'd156;
Cp[26] <= 11'd1010; Sp[26] <= 11'd162;
Cp[27] <= 11'd1009; Sp[27] <= 11'd169;
Cp[28] <= 11'd1008; Sp[28] <= 11'd175;
Cp[29] <= 11'd1007; Sp[29] <= 11'd181;
Cp[30] <= 11'd1006; Sp[30] <= 11'd187;
Cp[31] <= 11'd1005; Sp[31] <= 11'd193;
Cp[32] <= 11'd1004; Sp[32] <= 11'd199;
Cp[33] <= 11'd1003; Sp[33] <= 11'd206;
Cp[34] <= 11'd1001; Sp[34] <= 11'd212;
Cp[35] <= 11'd1000; Sp[35] <= 11'd218;
Cp[36] <= 11'd999; Sp[36] <= 11'd224;
Cp[37] <= 11'd997; Sp[37] <= 11'd230;
Cp[38] <= 11'd996; Sp[38] <= 11'd236;
Cp[39] <= 11'd994; Sp[39] <= 11'd242;
Cp[40] <= 11'd993; Sp[40] <= 11'd249;
Cp[41] <= 11'd991; Sp[41] <= 11'd255;
Cp[42] <= 11'd990; Sp[42] <= 11'd261;
Cp[43] <= 11'd988; Sp[43] <= 11'd267;
Cp[44] <= 11'd986; Sp[44] <= 11'd273;
Cp[45] <= 11'd985; Sp[45] <= 11'd279;
Cp[46] <= 11'd983; Sp[46] <= 11'd285;
Cp[47] <= 11'd981; Sp[47] <= 11'd291;
Cp[48] <= 11'd979; Sp[48] <= 11'd297;
Cp[49] <= 11'd977; Sp[49] <= 11'd303;
Cp[50] <= 11'd976; Sp[50] <= 11'd309;
Cp[51] <= 11'd974; Sp[51] <= 11'd315;
Cp[52] <= 11'd972; Sp[52] <= 11'd321;
Cp[53] <= 11'd970; Sp[53] <= 11'd327;
Cp[54] <= 11'd968; Sp[54] <= 11'd333;
Cp[55] <= 11'd966; Sp[55] <= 11'd339;
Cp[56] <= 11'd964; Sp[56] <= 11'd345;
Cp[57] <= 11'd961; Sp[57] <= 11'd351;
Cp[58] <= 11'd959; Sp[58] <= 11'd357;
Cp[59] <= 11'd957; Sp[59] <= 11'd363;
Cp[60] <= 11'd955; Sp[60] <= 11'd368;
Cp[61] <= 11'd952; Sp[61] <= 11'd374;
Cp[62] <= 11'd950; Sp[62] <= 11'd380;
Cp[63] <= 11'd948; Sp[63] <= 11'd386;
Cp[64] <= 11'd945; Sp[64] <= 11'd392;
Cp[65] <= 11'd943; Sp[65] <= 11'd398;
Cp[66] <= 11'd941; Sp[66] <= 11'd403;
Cp[67] <= 11'd938; Sp[67] <= 11'd409;
Cp[68] <= 11'd935; Sp[68] <= 11'd415;
Cp[69] <= 11'd933; Sp[69] <= 11'd421;
Cp[70] <= 11'd930; Sp[70] <= 11'd426;
Cp[71] <= 11'd928; Sp[71] <= 11'd432;
Cp[72] <= 11'd925; Sp[72] <= 11'd438;
Cp[73] <= 11'd922; Sp[73] <= 11'd443;
Cp[74] <= 11'd920; Sp[74] <= 11'd449;
Cp[75] <= 11'd917; Sp[75] <= 11'd455;
Cp[76] <= 11'd914; Sp[76] <= 11'd460;
Cp[77] <= 11'd911; Sp[77] <= 11'd466;
Cp[78] <= 11'd908; Sp[78] <= 11'd472;
Cp[79] <= 11'd905; Sp[79] <= 11'd477;
Cp[80] <= 11'd902; Sp[80] <= 11'd483;
Cp[81] <= 11'd899; Sp[81] <= 11'd488;
Cp[82] <= 11'd896; Sp[82] <= 11'd494;
Cp[83] <= 11'd893; Sp[83] <= 11'd499;
Cp[84] <= 11'd890; Sp[84] <= 11'd505;
Cp[85] <= 11'd887; Sp[85] <= 11'd510;
Cp[86] <= 11'd884; Sp[86] <= 11'd516;
Cp[87] <= 11'd881; Sp[87] <= 11'd521;
Cp[88] <= 11'd878; Sp[88] <= 11'd526;
Cp[89] <= 11'd874; Sp[89] <= 11'd532;
Cp[90] <= 11'd871; Sp[90] <= 11'd537;
Cp[91] <= 11'd868; Sp[91] <= 11'd542;
Cp[92] <= 11'd864; Sp[92] <= 11'd548;
Cp[93] <= 11'd861; Sp[93] <= 11'd553;
Cp[94] <= 11'd858; Sp[94] <= 11'd558;
Cp[95] <= 11'd854; Sp[95] <= 11'd564;
Cp[96] <= 11'd851; Sp[96] <= 11'd569;
Cp[97] <= 11'd847; Sp[97] <= 11'd574;
Cp[98] <= 11'd844; Sp[98] <= 11'd579;
Cp[99] <= 11'd840; Sp[99] <= 11'd584;
Cp[100] <= 11'd836; Sp[100] <= 11'd590;
Cp[101] <= 11'd833; Sp[101] <= 11'd595;
Cp[102] <= 11'd829; Sp[102] <= 11'd600;
Cp[103] <= 11'd825; Sp[103] <= 11'd605;
Cp[104] <= 11'd822; Sp[104] <= 11'd610;
Cp[105] <= 11'd818; Sp[105] <= 11'd615;
Cp[106] <= 11'd814; Sp[106] <= 11'd620;
Cp[107] <= 11'd810; Sp[107] <= 11'd625;
Cp[108] <= 11'd806; Sp[108] <= 11'd630;
Cp[109] <= 11'd802; Sp[109] <= 11'd635;
Cp[110] <= 11'd799; Sp[110] <= 11'd640;
Cp[111] <= 11'd795; Sp[111] <= 11'd645;
Cp[112] <= 11'd791; Sp[112] <= 11'd650;
Cp[113] <= 11'd787; Sp[113] <= 11'd654;
Cp[114] <= 11'd783; Sp[114] <= 11'd659;
Cp[115] <= 11'd779; Sp[115] <= 11'd664;
Cp[116] <= 11'd774; Sp[116] <= 11'd669;
Cp[117] <= 11'd770; Sp[117] <= 11'd674;
Cp[118] <= 11'd766; Sp[118] <= 11'd678;
Cp[119] <= 11'd762; Sp[119] <= 11'd683;
Cp[120] <= 11'd758; Sp[120] <= 11'd688;
Cp[121] <= 11'd753; Sp[121] <= 11'd692;
Cp[122] <= 11'd749; Sp[122] <= 11'd697;
Cp[123] <= 11'd745; Sp[123] <= 11'd702;
Cp[124] <= 11'd741; Sp[124] <= 11'd706;
Cp[125] <= 11'd736; Sp[125] <= 11'd711;
Cp[126] <= 11'd732; Sp[126] <= 11'd715;
Cp[127] <= 11'd727; Sp[127] <= 11'd720;
Cp[128] <= 11'd723; Sp[128] <= 11'd724;
Cp[129] <= 11'd719; Sp[129] <= 11'd729;
Cp[130] <= 11'd714; Sp[130] <= 11'd733;
Cp[131] <= 11'd710; Sp[131] <= 11'd737;
Cp[132] <= 11'd705; Sp[132] <= 11'd742;
Cp[133] <= 11'd700; Sp[133] <= 11'd746;
Cp[134] <= 11'd696; Sp[134] <= 11'd750;
Cp[135] <= 11'd691; Sp[135] <= 11'd755;
Cp[136] <= 11'd687; Sp[136] <= 11'd759;
Cp[137] <= 11'd682; Sp[137] <= 11'd763;
Cp[138] <= 11'd677; Sp[138] <= 11'd767;
Cp[139] <= 11'd672; Sp[139] <= 11'd771;
Cp[140] <= 11'd668; Sp[140] <= 11'd775;
Cp[141] <= 11'd663; Sp[141] <= 11'd780;
Cp[142] <= 11'd658; Sp[142] <= 11'd784;
Cp[143] <= 11'd653; Sp[143] <= 11'd788;
Cp[144] <= 11'd648; Sp[144] <= 11'd792;
Cp[145] <= 11'd644; Sp[145] <= 11'd796;
Cp[146] <= 11'd639; Sp[146] <= 11'd800;
Cp[147] <= 11'd634; Sp[147] <= 11'd803;
Cp[148] <= 11'd629; Sp[148] <= 11'd807;
Cp[149] <= 11'd624; Sp[149] <= 11'd811;
Cp[150] <= 11'd619; Sp[150] <= 11'd815;
Cp[151] <= 11'd614; Sp[151] <= 11'd819;
Cp[152] <= 11'd609; Sp[152] <= 11'd823;
Cp[153] <= 11'd604; Sp[153] <= 11'd826;
Cp[154] <= 11'd599; Sp[154] <= 11'd830;
Cp[155] <= 11'd593; Sp[155] <= 11'd834;
Cp[156] <= 11'd588; Sp[156] <= 11'd837;
Cp[157] <= 11'd583; Sp[157] <= 11'd841;
Cp[158] <= 11'd578; Sp[158] <= 11'd844;
Cp[159] <= 11'd573; Sp[159] <= 11'd848;
Cp[160] <= 11'd568; Sp[160] <= 11'd851;
Cp[161] <= 11'd562; Sp[161] <= 11'd855;
Cp[162] <= 11'd557; Sp[162] <= 11'd858;
Cp[163] <= 11'd552; Sp[163] <= 11'd862;
Cp[164] <= 11'd546; Sp[164] <= 11'd865;
Cp[165] <= 11'd541; Sp[165] <= 11'd869;
Cp[166] <= 11'd536; Sp[166] <= 11'd872;
Cp[167] <= 11'd530; Sp[167] <= 11'd875;
Cp[168] <= 11'd525; Sp[168] <= 11'd878;
Cp[169] <= 11'd520; Sp[169] <= 11'd882;
Cp[170] <= 11'd514; Sp[170] <= 11'd885;
Cp[171] <= 11'd509; Sp[171] <= 11'd888;
Cp[172] <= 11'd503; Sp[172] <= 11'd891;
Cp[173] <= 11'd498; Sp[173] <= 11'd894;
Cp[174] <= 11'd492; Sp[174] <= 11'd897;
Cp[175] <= 11'd487; Sp[175] <= 11'd900;
Cp[176] <= 11'd481; Sp[176] <= 11'd903;
Cp[177] <= 11'd476; Sp[177] <= 11'd906;
Cp[178] <= 11'd470; Sp[178] <= 11'd909;
Cp[179] <= 11'd465; Sp[179] <= 11'd912;
Cp[180] <= 11'd459; Sp[180] <= 11'd915;
Cp[181] <= 11'd453; Sp[181] <= 11'd917;
Cp[182] <= 11'd448; Sp[182] <= 11'd920;
Cp[183] <= 11'd442; Sp[183] <= 11'd923;
Cp[184] <= 11'd436; Sp[184] <= 11'd926;
Cp[185] <= 11'd431; Sp[185] <= 11'd928;
Cp[186] <= 11'd425; Sp[186] <= 11'd931;
Cp[187] <= 11'd419; Sp[187] <= 11'd934;
Cp[188] <= 11'd413; Sp[188] <= 11'd936;
Cp[189] <= 11'd408; Sp[189] <= 11'd939;
Cp[190] <= 11'd402; Sp[190] <= 11'd941;
Cp[191] <= 11'd396; Sp[191] <= 11'd944;
Cp[192] <= 11'd390; Sp[192] <= 11'd946;
Cp[193] <= 11'd384; Sp[193] <= 11'd948;
Cp[194] <= 11'd379; Sp[194] <= 11'd951;
Cp[195] <= 11'd373; Sp[195] <= 11'd953;
Cp[196] <= 11'd367; Sp[196] <= 11'd955;
Cp[197] <= 11'd361; Sp[197] <= 11'd958;
Cp[198] <= 11'd355; Sp[198] <= 11'd960;
Cp[199] <= 11'd349; Sp[199] <= 11'd962;
Cp[200] <= 11'd343; Sp[200] <= 11'd964;
Cp[201] <= 11'd337; Sp[201] <= 11'd966;
Cp[202] <= 11'd331; Sp[202] <= 11'd968;
Cp[203] <= 11'd325; Sp[203] <= 11'd970;
Cp[204] <= 11'd320; Sp[204] <= 11'd972;
Cp[205] <= 11'd314; Sp[205] <= 11'd974;
Cp[206] <= 11'd308; Sp[206] <= 11'd976;
Cp[207] <= 11'd302; Sp[207] <= 11'd978;
Cp[208] <= 11'd296; Sp[208] <= 11'd980;
Cp[209] <= 11'd290; Sp[209] <= 11'd982;
Cp[210] <= 11'd283; Sp[210] <= 11'd983;
Cp[211] <= 11'd277; Sp[211] <= 11'd985;
Cp[212] <= 11'd271; Sp[212] <= 11'd987;
Cp[213] <= 11'd265; Sp[213] <= 11'd988;
Cp[214] <= 11'd259; Sp[214] <= 11'd990;
Cp[215] <= 11'd253; Sp[215] <= 11'd992;
Cp[216] <= 11'd247; Sp[216] <= 11'd993;
Cp[217] <= 11'd241; Sp[217] <= 11'd995;
Cp[218] <= 11'd235; Sp[218] <= 11'd996;
Cp[219] <= 11'd229; Sp[219] <= 11'd998;
Cp[220] <= 11'd223; Sp[220] <= 11'd999;
Cp[221] <= 11'd216; Sp[221] <= 11'd1000;
Cp[222] <= 11'd210; Sp[222] <= 11'd1002;
Cp[223] <= 11'd204; Sp[223] <= 11'd1003;
Cp[224] <= 11'd198; Sp[224] <= 11'd1004;
Cp[225] <= 11'd192; Sp[225] <= 11'd1005;
Cp[226] <= 11'd186; Sp[226] <= 11'd1006;
Cp[227] <= 11'd179; Sp[227] <= 11'd1008;
Cp[228] <= 11'd173; Sp[228] <= 11'd1009;
Cp[229] <= 11'd167; Sp[229] <= 11'd1010;
Cp[230] <= 11'd161; Sp[230] <= 11'd1011;
Cp[231] <= 11'd155; Sp[231] <= 11'd1012;
Cp[232] <= 11'd148; Sp[232] <= 11'd1013;
Cp[233] <= 11'd142; Sp[233] <= 11'd1014;
Cp[234] <= 11'd136; Sp[234] <= 11'd1014;
Cp[235] <= 11'd130; Sp[235] <= 11'd1015;
Cp[236] <= 11'd123; Sp[236] <= 11'd1016;
Cp[237] <= 11'd117; Sp[237] <= 11'd1017;
Cp[238] <= 11'd111; Sp[238] <= 11'd1017;
Cp[239] <= 11'd105; Sp[239] <= 11'd1018;
Cp[240] <= 11'd98; Sp[240] <= 11'd1019;
Cp[241] <= 11'd92; Sp[241] <= 11'd1019;
Cp[242] <= 11'd86; Sp[242] <= 11'd1020;
Cp[243] <= 11'd80; Sp[243] <= 11'd1020;
Cp[244] <= 11'd73; Sp[244] <= 11'd1021;
Cp[245] <= 11'd67; Sp[245] <= 11'd1021;
Cp[246] <= 11'd61; Sp[246] <= 11'd1022;
Cp[247] <= 11'd55; Sp[247] <= 11'd1022;
Cp[248] <= 11'd48; Sp[248] <= 11'd1022;
Cp[249] <= 11'd42; Sp[249] <= 11'd1023;
Cp[250] <= 11'd36; Sp[250] <= 11'd1023;
Cp[251] <= 11'd29; Sp[251] <= 11'd1023;
Cp[252] <= 11'd23; Sp[252] <= 11'd1023;
Cp[253] <= 11'd17; Sp[253] <= 11'd1023;
Cp[254] <= 11'd11; Sp[254] <= 11'd1023;
Cp[255] <= 11'd4; Sp[255] <= 11'd1023;
Cp[256] <= -11'd1; Sp[256] <= 11'd1023;
Cp[257] <= -11'd7; Sp[257] <= 11'd1023;
Cp[258] <= -11'd14; Sp[258] <= 11'd1023;
Cp[259] <= -11'd20; Sp[259] <= 11'd1023;
Cp[260] <= -11'd26; Sp[260] <= 11'd1023;
Cp[261] <= -11'd33; Sp[261] <= 11'd1023;
Cp[262] <= -11'd39; Sp[262] <= 11'd1023;
Cp[263] <= -11'd45; Sp[263] <= 11'd1022;
Cp[264] <= -11'd51; Sp[264] <= 11'd1022;
Cp[265] <= -11'd58; Sp[265] <= 11'd1022;
Cp[266] <= -11'd64; Sp[266] <= 11'd1021;
Cp[267] <= -11'd70; Sp[267] <= 11'd1021;
Cp[268] <= -11'd76; Sp[268] <= 11'd1021;
Cp[269] <= -11'd83; Sp[269] <= 11'd1020;
Cp[270] <= -11'd89; Sp[270] <= 11'd1020;
Cp[271] <= -11'd95; Sp[271] <= 11'd1019;
Cp[272] <= -11'd102; Sp[272] <= 11'd1018;
Cp[273] <= -11'd108; Sp[273] <= 11'd1018;
Cp[274] <= -11'd114; Sp[274] <= 11'd1017;
Cp[275] <= -11'd120; Sp[275] <= 11'd1016;
Cp[276] <= -11'd127; Sp[276] <= 11'd1016;
Cp[277] <= -11'd133; Sp[277] <= 11'd1015;
Cp[278] <= -11'd139; Sp[278] <= 11'd1014;
Cp[279] <= -11'd145; Sp[279] <= 11'd1013;
Cp[280] <= -11'd151; Sp[280] <= 11'd1012;
Cp[281] <= -11'd158; Sp[281] <= 11'd1011;
Cp[282] <= -11'd164; Sp[282] <= 11'd1010;
Cp[283] <= -11'd170; Sp[283] <= 11'd1009;
Cp[284] <= -11'd176; Sp[284] <= 11'd1008;
Cp[285] <= -11'd182; Sp[285] <= 11'd1007;
Cp[286] <= -11'd189; Sp[286] <= 11'd1006;
Cp[287] <= -11'd195; Sp[287] <= 11'd1005;
Cp[288] <= -11'd201; Sp[288] <= 11'd1003;
Cp[289] <= -11'd207; Sp[289] <= 11'd1002;
Cp[290] <= -11'd213; Sp[290] <= 11'd1001;
Cp[291] <= -11'd219; Sp[291] <= 11'd1000;
Cp[292] <= -11'd226; Sp[292] <= 11'd998;
Cp[293] <= -11'd232; Sp[293] <= 11'd997;
Cp[294] <= -11'd238; Sp[294] <= 11'd995;
Cp[295] <= -11'd244; Sp[295] <= 11'd994;
Cp[296] <= -11'd250; Sp[296] <= 11'd992;
Cp[297] <= -11'd256; Sp[297] <= 11'd991;
Cp[298] <= -11'd262; Sp[298] <= 11'd989;
Cp[299] <= -11'd268; Sp[299] <= 11'd988;
Cp[300] <= -11'd274; Sp[300] <= 11'd986;
Cp[301] <= -11'd280; Sp[301] <= 11'd984;
Cp[302] <= -11'd286; Sp[302] <= 11'd982;
Cp[303] <= -11'd293; Sp[303] <= 11'd981;
Cp[304] <= -11'd299; Sp[304] <= 11'd979;
Cp[305] <= -11'd305; Sp[305] <= 11'd977;
Cp[306] <= -11'd311; Sp[306] <= 11'd975;
Cp[307] <= -11'd317; Sp[307] <= 11'd973;
Cp[308] <= -11'd323; Sp[308] <= 11'd971;
Cp[309] <= -11'd328; Sp[309] <= 11'd969;
Cp[310] <= -11'd334; Sp[310] <= 11'd967;
Cp[311] <= -11'd340; Sp[311] <= 11'd965;
Cp[312] <= -11'd346; Sp[312] <= 11'd963;
Cp[313] <= -11'd352; Sp[313] <= 11'd961;
Cp[314] <= -11'd358; Sp[314] <= 11'd959;
Cp[315] <= -11'd364; Sp[315] <= 11'd956;
Cp[316] <= -11'd370; Sp[316] <= 11'd954;
Cp[317] <= -11'd376; Sp[317] <= 11'd952;
Cp[318] <= -11'd382; Sp[318] <= 11'd950;
Cp[319] <= -11'd387; Sp[319] <= 11'd947;
Cp[320] <= -11'd393; Sp[320] <= 11'd945;
Cp[321] <= -11'd399; Sp[321] <= 11'd942;
Cp[322] <= -11'd405; Sp[322] <= 11'd940;
Cp[323] <= -11'd411; Sp[323] <= 11'd937;
Cp[324] <= -11'd416; Sp[324] <= 11'd935;
Cp[325] <= -11'd422; Sp[325] <= 11'd932;
Cp[326] <= -11'd428; Sp[326] <= 11'd930;
Cp[327] <= -11'd433; Sp[327] <= 11'd927;
Cp[328] <= -11'd439; Sp[328] <= 11'd924;
Cp[329] <= -11'd445; Sp[329] <= 11'd922;
Cp[330] <= -11'd450; Sp[330] <= 11'd919;
Cp[331] <= -11'd456; Sp[331] <= 11'd916;
Cp[332] <= -11'd462; Sp[332] <= 11'd913;
Cp[333] <= -11'd467; Sp[333] <= 11'd910;
Cp[334] <= -11'd473; Sp[334] <= 11'd907;
Cp[335] <= -11'd478; Sp[335] <= 11'd905;
Cp[336] <= -11'd484; Sp[336] <= 11'd902;
Cp[337] <= -11'd490; Sp[337] <= 11'd899;
Cp[338] <= -11'd495; Sp[338] <= 11'd896;
Cp[339] <= -11'd501; Sp[339] <= 11'd893;
Cp[340] <= -11'd506; Sp[340] <= 11'd889;
Cp[341] <= -11'd511; Sp[341] <= 11'd886;
Cp[342] <= -11'd517; Sp[342] <= 11'd883;
Cp[343] <= -11'd522; Sp[343] <= 11'd880;
Cp[344] <= -11'd528; Sp[344] <= 11'd877;
Cp[345] <= -11'd533; Sp[345] <= 11'd873;
Cp[346] <= -11'd538; Sp[346] <= 11'd870;
Cp[347] <= -11'd544; Sp[347] <= 11'd867;
Cp[348] <= -11'd549; Sp[348] <= 11'd863;
Cp[349] <= -11'd554; Sp[349] <= 11'd860;
Cp[350] <= -11'd560; Sp[350] <= 11'd857;
Cp[351] <= -11'd565; Sp[351] <= 11'd853;
Cp[352] <= -11'd570; Sp[352] <= 11'd850;
Cp[353] <= -11'd575; Sp[353] <= 11'd846;
Cp[354] <= -11'd581; Sp[354] <= 11'd843;
Cp[355] <= -11'd586; Sp[355] <= 11'd839;
Cp[356] <= -11'd591; Sp[356] <= 11'd835;
Cp[357] <= -11'd596; Sp[357] <= 11'd832;
Cp[358] <= -11'd601; Sp[358] <= 11'd828;
Cp[359] <= -11'd606; Sp[359] <= 11'd824;
Cp[360] <= -11'd611; Sp[360] <= 11'd821;
Cp[361] <= -11'd616; Sp[361] <= 11'd817;
Cp[362] <= -11'd621; Sp[362] <= 11'd813;
Cp[363] <= -11'd626; Sp[363] <= 11'd809;
Cp[364] <= -11'd631; Sp[364] <= 11'd805;
Cp[365] <= -11'd636; Sp[365] <= 11'd801;
Cp[366] <= -11'd641; Sp[366] <= 11'd798;
Cp[367] <= -11'd646; Sp[367] <= 11'd794;
Cp[368] <= -11'd651; Sp[368] <= 11'd790;
Cp[369] <= -11'd656; Sp[369] <= 11'd786;
Cp[370] <= -11'd661; Sp[370] <= 11'd782;
Cp[371] <= -11'd665; Sp[371] <= 11'd777;
Cp[372] <= -11'd670; Sp[372] <= 11'd773;
Cp[373] <= -11'd675; Sp[373] <= 11'd769;
Cp[374] <= -11'd680; Sp[374] <= 11'd765;
Cp[375] <= -11'd684; Sp[375] <= 11'd761;
Cp[376] <= -11'd689; Sp[376] <= 11'd757;
Cp[377] <= -11'd694; Sp[377] <= 11'd752;
Cp[378] <= -11'd698; Sp[378] <= 11'd748;
Cp[379] <= -11'd703; Sp[379] <= 11'd744;
Cp[380] <= -11'd707; Sp[380] <= 11'd740;
Cp[381] <= -11'd712; Sp[381] <= 11'd735;
Cp[382] <= -11'd716; Sp[382] <= 11'd731;
Cp[383] <= -11'd721; Sp[383] <= 11'd726;
Cp[384] <= -11'd725; Sp[384] <= 11'd722;
Cp[385] <= -11'd730; Sp[385] <= 11'd717;
Cp[386] <= -11'd734; Sp[386] <= 11'd713;
Cp[387] <= -11'd738; Sp[387] <= 11'd708;
Cp[388] <= -11'd743; Sp[388] <= 11'd704;
Cp[389] <= -11'd747; Sp[389] <= 11'd699;
Cp[390] <= -11'd751; Sp[390] <= 11'd695;
Cp[391] <= -11'd756; Sp[391] <= 11'd690;
Cp[392] <= -11'd760; Sp[392] <= 11'd685;
Cp[393] <= -11'd764; Sp[393] <= 11'd681;
Cp[394] <= -11'd768; Sp[394] <= 11'd676;
Cp[395] <= -11'd772; Sp[395] <= 11'd671;
Cp[396] <= -11'd776; Sp[396] <= 11'd667;
Cp[397] <= -11'd781; Sp[397] <= 11'd662;
Cp[398] <= -11'd785; Sp[398] <= 11'd657;
Cp[399] <= -11'd789; Sp[399] <= 11'd652;
Cp[400] <= -11'd793; Sp[400] <= 11'd647;
Cp[401] <= -11'd797; Sp[401] <= 11'd642;
Cp[402] <= -11'd801; Sp[402] <= 11'd637;
Cp[403] <= -11'd804; Sp[403] <= 11'd632;
Cp[404] <= -11'd808; Sp[404] <= 11'd628;
Cp[405] <= -11'd812; Sp[405] <= 11'd623;
Cp[406] <= -11'd816; Sp[406] <= 11'd618;
Cp[407] <= -11'd820; Sp[407] <= 11'd613;
Cp[408] <= -11'd823; Sp[408] <= 11'd607;
Cp[409] <= -11'd827; Sp[409] <= 11'd602;
Cp[410] <= -11'd831; Sp[410] <= 11'd597;
Cp[411] <= -11'd835; Sp[411] <= 11'd592;
Cp[412] <= -11'd838; Sp[412] <= 11'd587;
Cp[413] <= -11'd842; Sp[413] <= 11'd582;
Cp[414] <= -11'd845; Sp[414] <= 11'd577;
Cp[415] <= -11'd849; Sp[415] <= 11'd572;
Cp[416] <= -11'd852; Sp[416] <= 11'd566;
Cp[417] <= -11'd856; Sp[417] <= 11'd561;
Cp[418] <= -11'd859; Sp[418] <= 11'd556;
Cp[419] <= -11'd863; Sp[419] <= 11'd550;
Cp[420] <= -11'd866; Sp[420] <= 11'd545;
Cp[421] <= -11'd869; Sp[421] <= 11'd540;
Cp[422] <= -11'd873; Sp[422] <= 11'd534;
Cp[423] <= -11'd876; Sp[423] <= 11'd529;
Cp[424] <= -11'd879; Sp[424] <= 11'd524;
Cp[425] <= -11'd882; Sp[425] <= 11'd518;
Cp[426] <= -11'd886; Sp[426] <= 11'd513;
Cp[427] <= -11'd889; Sp[427] <= 11'd507;
Cp[428] <= -11'd892; Sp[428] <= 11'd502;
Cp[429] <= -11'd895; Sp[429] <= 11'd496;
Cp[430] <= -11'd898; Sp[430] <= 11'd491;
Cp[431] <= -11'd901; Sp[431] <= 11'd485;
Cp[432] <= -11'd904; Sp[432] <= 11'd480;
Cp[433] <= -11'd907; Sp[433] <= 11'd474;
Cp[434] <= -11'd910; Sp[434] <= 11'd469;
Cp[435] <= -11'd913; Sp[435] <= 11'd463;
Cp[436] <= -11'd915; Sp[436] <= 11'd458;
Cp[437] <= -11'd918; Sp[437] <= 11'd452;
Cp[438] <= -11'd921; Sp[438] <= 11'd446;
Cp[439] <= -11'd924; Sp[439] <= 11'd441;
Cp[440] <= -11'd926; Sp[440] <= 11'd435;
Cp[441] <= -11'd929; Sp[441] <= 11'd429;
Cp[442] <= -11'd932; Sp[442] <= 11'd423;
Cp[443] <= -11'd934; Sp[443] <= 11'd418;
Cp[444] <= -11'd937; Sp[444] <= 11'd412;
Cp[445] <= -11'd939; Sp[445] <= 11'd406;
Cp[446] <= -11'd942; Sp[446] <= 11'd400;
Cp[447] <= -11'd944; Sp[447] <= 11'd395;
Cp[448] <= -11'd947; Sp[448] <= 11'd389;
Cp[449] <= -11'd949; Sp[449] <= 11'd383;
Cp[450] <= -11'd951; Sp[450] <= 11'd377;
Cp[451] <= -11'd954; Sp[451] <= 11'd371;
Cp[452] <= -11'd956; Sp[452] <= 11'd365;
Cp[453] <= -11'd958; Sp[453] <= 11'd360;
Cp[454] <= -11'd960; Sp[454] <= 11'd354;
Cp[455] <= -11'd962; Sp[455] <= 11'd348;
Cp[456] <= -11'd965; Sp[456] <= 11'd342;
Cp[457] <= -11'd967; Sp[457] <= 11'd336;
Cp[458] <= -11'd969; Sp[458] <= 11'd330;
Cp[459] <= -11'd971; Sp[459] <= 11'd324;
Cp[460] <= -11'd973; Sp[460] <= 11'd318;
Cp[461] <= -11'd975; Sp[461] <= 11'd312;
Cp[462] <= -11'd977; Sp[462] <= 11'd306;
Cp[463] <= -11'd978; Sp[463] <= 11'd300;
Cp[464] <= -11'd980; Sp[464] <= 11'd294;
Cp[465] <= -11'd982; Sp[465] <= 11'd288;
Cp[466] <= -11'd984; Sp[466] <= 11'd282;
Cp[467] <= -11'd985; Sp[467] <= 11'd276;
Cp[468] <= -11'd987; Sp[468] <= 11'd270;
Cp[469] <= -11'd989; Sp[469] <= 11'd264;
Cp[470] <= -11'd990; Sp[470] <= 11'd258;
Cp[471] <= -11'd992; Sp[471] <= 11'd252;
Cp[472] <= -11'd994; Sp[472] <= 11'd245;
Cp[473] <= -11'd995; Sp[473] <= 11'd239;
Cp[474] <= -11'd996; Sp[474] <= 11'd233;
Cp[475] <= -11'd998; Sp[475] <= 11'd227;
Cp[476] <= -11'd999; Sp[476] <= 11'd221;
Cp[477] <= -11'd1001; Sp[477] <= 11'd215;
Cp[478] <= -11'd1002; Sp[478] <= 11'd209;
Cp[479] <= -11'd1003; Sp[479] <= 11'd203;
Cp[480] <= -11'd1004; Sp[480] <= 11'd196;
Cp[481] <= -11'd1006; Sp[481] <= 11'd190;
Cp[482] <= -11'd1007; Sp[482] <= 11'd184;
Cp[483] <= -11'd1008; Sp[483] <= 11'd178;
Cp[484] <= -11'd1009; Sp[484] <= 11'd172;
Cp[485] <= -11'd1010; Sp[485] <= 11'd165;
Cp[486] <= -11'd1011; Sp[486] <= 11'd159;
Cp[487] <= -11'd1012; Sp[487] <= 11'd153;
Cp[488] <= -11'd1013; Sp[488] <= 11'd147;
Cp[489] <= -11'd1014; Sp[489] <= 11'd141;
Cp[490] <= -11'd1015; Sp[490] <= 11'd134;
Cp[491] <= -11'd1015; Sp[491] <= 11'd128;
Cp[492] <= -11'd1016; Sp[492] <= 11'd122;
Cp[493] <= -11'd1017; Sp[493] <= 11'd116;
Cp[494] <= -11'd1018; Sp[494] <= 11'd109;
Cp[495] <= -11'd1018; Sp[495] <= 11'd103;
Cp[496] <= -11'd1019; Sp[496] <= 11'd97;
Cp[497] <= -11'd1019; Sp[497] <= 11'd91;
Cp[498] <= -11'd1020; Sp[498] <= 11'd84;
Cp[499] <= -11'd1020; Sp[499] <= 11'd78;
Cp[500] <= -11'd1021; Sp[500] <= 11'd72;
Cp[501] <= -11'd1021; Sp[501] <= 11'd65;
Cp[502] <= -11'd1022; Sp[502] <= 11'd59;
Cp[503] <= -11'd1022; Sp[503] <= 11'd53;
Cp[504] <= -11'd1022; Sp[504] <= 11'd47;
Cp[505] <= -11'd1023; Sp[505] <= 11'd40;
Cp[506] <= -11'd1023; Sp[506] <= 11'd34;
Cp[507] <= -11'd1023; Sp[507] <= 11'd28;
Cp[508] <= -11'd1023; Sp[508] <= 11'd22;
Cp[509] <= -11'd1023; Sp[509] <= 11'd15;
Cp[510] <= -11'd1023; Sp[510] <= 11'd9;
Cp[511] <= -11'd1023; Sp[511] <= 11'd3;
Cp[512] <= -11'd1023; Sp[512] <= -11'd3;
Cp[513] <= -11'd1023; Sp[513] <= -11'd9;
Cp[514] <= -11'd1023; Sp[514] <= -11'd15;
Cp[515] <= -11'd1023; Sp[515] <= -11'd22;
Cp[516] <= -11'd1023; Sp[516] <= -11'd28;
Cp[517] <= -11'd1023; Sp[517] <= -11'd34;
Cp[518] <= -11'd1023; Sp[518] <= -11'd40;
Cp[519] <= -11'd1022; Sp[519] <= -11'd47;
Cp[520] <= -11'd1022; Sp[520] <= -11'd53;
Cp[521] <= -11'd1022; Sp[521] <= -11'd59;
Cp[522] <= -11'd1021; Sp[522] <= -11'd65;
Cp[523] <= -11'd1021; Sp[523] <= -11'd72;
Cp[524] <= -11'd1020; Sp[524] <= -11'd78;
Cp[525] <= -11'd1020; Sp[525] <= -11'd84;
Cp[526] <= -11'd1019; Sp[526] <= -11'd91;
Cp[527] <= -11'd1019; Sp[527] <= -11'd97;
Cp[528] <= -11'd1018; Sp[528] <= -11'd103;
Cp[529] <= -11'd1018; Sp[529] <= -11'd109;
Cp[530] <= -11'd1017; Sp[530] <= -11'd116;
Cp[531] <= -11'd1016; Sp[531] <= -11'd122;
Cp[532] <= -11'd1015; Sp[532] <= -11'd128;
Cp[533] <= -11'd1015; Sp[533] <= -11'd134;
Cp[534] <= -11'd1014; Sp[534] <= -11'd141;
Cp[535] <= -11'd1013; Sp[535] <= -11'd147;
Cp[536] <= -11'd1012; Sp[536] <= -11'd153;
Cp[537] <= -11'd1011; Sp[537] <= -11'd159;
Cp[538] <= -11'd1010; Sp[538] <= -11'd165;
Cp[539] <= -11'd1009; Sp[539] <= -11'd172;
Cp[540] <= -11'd1008; Sp[540] <= -11'd178;
Cp[541] <= -11'd1007; Sp[541] <= -11'd184;
Cp[542] <= -11'd1006; Sp[542] <= -11'd190;
Cp[543] <= -11'd1004; Sp[543] <= -11'd196;
Cp[544] <= -11'd1003; Sp[544] <= -11'd203;
Cp[545] <= -11'd1002; Sp[545] <= -11'd209;
Cp[546] <= -11'd1001; Sp[546] <= -11'd215;
Cp[547] <= -11'd999; Sp[547] <= -11'd221;
Cp[548] <= -11'd998; Sp[548] <= -11'd227;
Cp[549] <= -11'd996; Sp[549] <= -11'd233;
Cp[550] <= -11'd995; Sp[550] <= -11'd239;
Cp[551] <= -11'd994; Sp[551] <= -11'd245;
Cp[552] <= -11'd992; Sp[552] <= -11'd252;
Cp[553] <= -11'd990; Sp[553] <= -11'd258;
Cp[554] <= -11'd989; Sp[554] <= -11'd264;
Cp[555] <= -11'd987; Sp[555] <= -11'd270;
Cp[556] <= -11'd985; Sp[556] <= -11'd276;
Cp[557] <= -11'd984; Sp[557] <= -11'd282;
Cp[558] <= -11'd982; Sp[558] <= -11'd288;
Cp[559] <= -11'd980; Sp[559] <= -11'd294;
Cp[560] <= -11'd978; Sp[560] <= -11'd300;
Cp[561] <= -11'd977; Sp[561] <= -11'd306;
Cp[562] <= -11'd975; Sp[562] <= -11'd312;
Cp[563] <= -11'd973; Sp[563] <= -11'd318;
Cp[564] <= -11'd971; Sp[564] <= -11'd324;
Cp[565] <= -11'd969; Sp[565] <= -11'd330;
Cp[566] <= -11'd967; Sp[566] <= -11'd336;
Cp[567] <= -11'd965; Sp[567] <= -11'd342;
Cp[568] <= -11'd962; Sp[568] <= -11'd348;
Cp[569] <= -11'd960; Sp[569] <= -11'd354;
Cp[570] <= -11'd958; Sp[570] <= -11'd360;
Cp[571] <= -11'd956; Sp[571] <= -11'd365;
Cp[572] <= -11'd954; Sp[572] <= -11'd371;
Cp[573] <= -11'd951; Sp[573] <= -11'd377;
Cp[574] <= -11'd949; Sp[574] <= -11'd383;
Cp[575] <= -11'd947; Sp[575] <= -11'd389;
Cp[576] <= -11'd944; Sp[576] <= -11'd395;
Cp[577] <= -11'd942; Sp[577] <= -11'd400;
Cp[578] <= -11'd939; Sp[578] <= -11'd406;
Cp[579] <= -11'd937; Sp[579] <= -11'd412;
Cp[580] <= -11'd934; Sp[580] <= -11'd418;
Cp[581] <= -11'd932; Sp[581] <= -11'd423;
Cp[582] <= -11'd929; Sp[582] <= -11'd429;
Cp[583] <= -11'd926; Sp[583] <= -11'd435;
Cp[584] <= -11'd924; Sp[584] <= -11'd441;
Cp[585] <= -11'd921; Sp[585] <= -11'd446;
Cp[586] <= -11'd918; Sp[586] <= -11'd452;
Cp[587] <= -11'd915; Sp[587] <= -11'd458;
Cp[588] <= -11'd913; Sp[588] <= -11'd463;
Cp[589] <= -11'd910; Sp[589] <= -11'd469;
Cp[590] <= -11'd907; Sp[590] <= -11'd474;
Cp[591] <= -11'd904; Sp[591] <= -11'd480;
Cp[592] <= -11'd901; Sp[592] <= -11'd485;
Cp[593] <= -11'd898; Sp[593] <= -11'd491;
Cp[594] <= -11'd895; Sp[594] <= -11'd496;
Cp[595] <= -11'd892; Sp[595] <= -11'd502;
Cp[596] <= -11'd889; Sp[596] <= -11'd507;
Cp[597] <= -11'd886; Sp[597] <= -11'd513;
Cp[598] <= -11'd882; Sp[598] <= -11'd518;
Cp[599] <= -11'd879; Sp[599] <= -11'd524;
Cp[600] <= -11'd876; Sp[600] <= -11'd529;
Cp[601] <= -11'd873; Sp[601] <= -11'd534;
Cp[602] <= -11'd869; Sp[602] <= -11'd540;
Cp[603] <= -11'd866; Sp[603] <= -11'd545;
Cp[604] <= -11'd863; Sp[604] <= -11'd550;
Cp[605] <= -11'd859; Sp[605] <= -11'd556;
Cp[606] <= -11'd856; Sp[606] <= -11'd561;
Cp[607] <= -11'd852; Sp[607] <= -11'd566;
Cp[608] <= -11'd849; Sp[608] <= -11'd572;
Cp[609] <= -11'd845; Sp[609] <= -11'd577;
Cp[610] <= -11'd842; Sp[610] <= -11'd582;
Cp[611] <= -11'd838; Sp[611] <= -11'd587;
Cp[612] <= -11'd835; Sp[612] <= -11'd592;
Cp[613] <= -11'd831; Sp[613] <= -11'd597;
Cp[614] <= -11'd827; Sp[614] <= -11'd602;
Cp[615] <= -11'd823; Sp[615] <= -11'd607;
Cp[616] <= -11'd820; Sp[616] <= -11'd613;
Cp[617] <= -11'd816; Sp[617] <= -11'd618;
Cp[618] <= -11'd812; Sp[618] <= -11'd623;
Cp[619] <= -11'd808; Sp[619] <= -11'd628;
Cp[620] <= -11'd804; Sp[620] <= -11'd632;
Cp[621] <= -11'd801; Sp[621] <= -11'd637;
Cp[622] <= -11'd797; Sp[622] <= -11'd642;
Cp[623] <= -11'd793; Sp[623] <= -11'd647;
Cp[624] <= -11'd789; Sp[624] <= -11'd652;
Cp[625] <= -11'd785; Sp[625] <= -11'd657;
Cp[626] <= -11'd781; Sp[626] <= -11'd662;
Cp[627] <= -11'd776; Sp[627] <= -11'd667;
Cp[628] <= -11'd772; Sp[628] <= -11'd671;
Cp[629] <= -11'd768; Sp[629] <= -11'd676;
Cp[630] <= -11'd764; Sp[630] <= -11'd681;
Cp[631] <= -11'd760; Sp[631] <= -11'd685;
Cp[632] <= -11'd756; Sp[632] <= -11'd690;
Cp[633] <= -11'd751; Sp[633] <= -11'd695;
Cp[634] <= -11'd747; Sp[634] <= -11'd699;
Cp[635] <= -11'd743; Sp[635] <= -11'd704;
Cp[636] <= -11'd738; Sp[636] <= -11'd708;
Cp[637] <= -11'd734; Sp[637] <= -11'd713;
Cp[638] <= -11'd730; Sp[638] <= -11'd717;
Cp[639] <= -11'd725; Sp[639] <= -11'd722;
Cp[640] <= -11'd721; Sp[640] <= -11'd726;
Cp[641] <= -11'd716; Sp[641] <= -11'd731;
Cp[642] <= -11'd712; Sp[642] <= -11'd735;
Cp[643] <= -11'd707; Sp[643] <= -11'd740;
Cp[644] <= -11'd703; Sp[644] <= -11'd744;
Cp[645] <= -11'd698; Sp[645] <= -11'd748;
Cp[646] <= -11'd694; Sp[646] <= -11'd752;
Cp[647] <= -11'd689; Sp[647] <= -11'd757;
Cp[648] <= -11'd684; Sp[648] <= -11'd761;
Cp[649] <= -11'd680; Sp[649] <= -11'd765;
Cp[650] <= -11'd675; Sp[650] <= -11'd769;
Cp[651] <= -11'd670; Sp[651] <= -11'd773;
Cp[652] <= -11'd665; Sp[652] <= -11'd777;
Cp[653] <= -11'd661; Sp[653] <= -11'd782;
Cp[654] <= -11'd656; Sp[654] <= -11'd786;
Cp[655] <= -11'd651; Sp[655] <= -11'd790;
Cp[656] <= -11'd646; Sp[656] <= -11'd794;
Cp[657] <= -11'd641; Sp[657] <= -11'd798;
Cp[658] <= -11'd636; Sp[658] <= -11'd801;
Cp[659] <= -11'd631; Sp[659] <= -11'd805;
Cp[660] <= -11'd626; Sp[660] <= -11'd809;
Cp[661] <= -11'd621; Sp[661] <= -11'd813;
Cp[662] <= -11'd616; Sp[662] <= -11'd817;
Cp[663] <= -11'd611; Sp[663] <= -11'd821;
Cp[664] <= -11'd606; Sp[664] <= -11'd824;
Cp[665] <= -11'd601; Sp[665] <= -11'd828;
Cp[666] <= -11'd596; Sp[666] <= -11'd832;
Cp[667] <= -11'd591; Sp[667] <= -11'd835;
Cp[668] <= -11'd586; Sp[668] <= -11'd839;
Cp[669] <= -11'd581; Sp[669] <= -11'd843;
Cp[670] <= -11'd575; Sp[670] <= -11'd846;
Cp[671] <= -11'd570; Sp[671] <= -11'd850;
Cp[672] <= -11'd565; Sp[672] <= -11'd853;
Cp[673] <= -11'd560; Sp[673] <= -11'd857;
Cp[674] <= -11'd554; Sp[674] <= -11'd860;
Cp[675] <= -11'd549; Sp[675] <= -11'd863;
Cp[676] <= -11'd544; Sp[676] <= -11'd867;
Cp[677] <= -11'd538; Sp[677] <= -11'd870;
Cp[678] <= -11'd533; Sp[678] <= -11'd873;
Cp[679] <= -11'd528; Sp[679] <= -11'd877;
Cp[680] <= -11'd522; Sp[680] <= -11'd880;
Cp[681] <= -11'd517; Sp[681] <= -11'd883;
Cp[682] <= -11'd512; Sp[682] <= -11'd886;
Cp[683] <= -11'd506; Sp[683] <= -11'd889;
Cp[684] <= -11'd501; Sp[684] <= -11'd893;
Cp[685] <= -11'd495; Sp[685] <= -11'd896;
Cp[686] <= -11'd490; Sp[686] <= -11'd899;
Cp[687] <= -11'd484; Sp[687] <= -11'd902;
Cp[688] <= -11'd478; Sp[688] <= -11'd905;
Cp[689] <= -11'd473; Sp[689] <= -11'd907;
Cp[690] <= -11'd467; Sp[690] <= -11'd910;
Cp[691] <= -11'd462; Sp[691] <= -11'd913;
Cp[692] <= -11'd456; Sp[692] <= -11'd916;
Cp[693] <= -11'd450; Sp[693] <= -11'd919;
Cp[694] <= -11'd445; Sp[694] <= -11'd922;
Cp[695] <= -11'd439; Sp[695] <= -11'd924;
Cp[696] <= -11'd433; Sp[696] <= -11'd927;
Cp[697] <= -11'd428; Sp[697] <= -11'd930;
Cp[698] <= -11'd422; Sp[698] <= -11'd932;
Cp[699] <= -11'd416; Sp[699] <= -11'd935;
Cp[700] <= -11'd411; Sp[700] <= -11'd937;
Cp[701] <= -11'd405; Sp[701] <= -11'd940;
Cp[702] <= -11'd399; Sp[702] <= -11'd942;
Cp[703] <= -11'd393; Sp[703] <= -11'd945;
Cp[704] <= -11'd387; Sp[704] <= -11'd947;
Cp[705] <= -11'd382; Sp[705] <= -11'd950;
Cp[706] <= -11'd376; Sp[706] <= -11'd952;
Cp[707] <= -11'd370; Sp[707] <= -11'd954;
Cp[708] <= -11'd364; Sp[708] <= -11'd956;
Cp[709] <= -11'd358; Sp[709] <= -11'd959;
Cp[710] <= -11'd352; Sp[710] <= -11'd961;
Cp[711] <= -11'd346; Sp[711] <= -11'd963;
Cp[712] <= -11'd340; Sp[712] <= -11'd965;
Cp[713] <= -11'd334; Sp[713] <= -11'd967;
Cp[714] <= -11'd328; Sp[714] <= -11'd969;
Cp[715] <= -11'd323; Sp[715] <= -11'd971;
Cp[716] <= -11'd317; Sp[716] <= -11'd973;
Cp[717] <= -11'd311; Sp[717] <= -11'd975;
Cp[718] <= -11'd305; Sp[718] <= -11'd977;
Cp[719] <= -11'd299; Sp[719] <= -11'd979;
Cp[720] <= -11'd293; Sp[720] <= -11'd981;
Cp[721] <= -11'd286; Sp[721] <= -11'd982;
Cp[722] <= -11'd280; Sp[722] <= -11'd984;
Cp[723] <= -11'd274; Sp[723] <= -11'd986;
Cp[724] <= -11'd268; Sp[724] <= -11'd988;
Cp[725] <= -11'd262; Sp[725] <= -11'd989;
Cp[726] <= -11'd256; Sp[726] <= -11'd991;
Cp[727] <= -11'd250; Sp[727] <= -11'd992;
Cp[728] <= -11'd244; Sp[728] <= -11'd994;
Cp[729] <= -11'd238; Sp[729] <= -11'd995;
Cp[730] <= -11'd232; Sp[730] <= -11'd997;
Cp[731] <= -11'd226; Sp[731] <= -11'd998;
Cp[732] <= -11'd219; Sp[732] <= -11'd1000;
Cp[733] <= -11'd213; Sp[733] <= -11'd1001;
Cp[734] <= -11'd207; Sp[734] <= -11'd1002;
Cp[735] <= -11'd201; Sp[735] <= -11'd1003;
Cp[736] <= -11'd195; Sp[736] <= -11'd1005;
Cp[737] <= -11'd189; Sp[737] <= -11'd1006;
Cp[738] <= -11'd182; Sp[738] <= -11'd1007;
Cp[739] <= -11'd176; Sp[739] <= -11'd1008;
Cp[740] <= -11'd170; Sp[740] <= -11'd1009;
Cp[741] <= -11'd164; Sp[741] <= -11'd1010;
Cp[742] <= -11'd158; Sp[742] <= -11'd1011;
Cp[743] <= -11'd151; Sp[743] <= -11'd1012;
Cp[744] <= -11'd145; Sp[744] <= -11'd1013;
Cp[745] <= -11'd139; Sp[745] <= -11'd1014;
Cp[746] <= -11'd133; Sp[746] <= -11'd1015;
Cp[747] <= -11'd127; Sp[747] <= -11'd1016;
Cp[748] <= -11'd120; Sp[748] <= -11'd1016;
Cp[749] <= -11'd114; Sp[749] <= -11'd1017;
Cp[750] <= -11'd108; Sp[750] <= -11'd1018;
Cp[751] <= -11'd102; Sp[751] <= -11'd1018;
Cp[752] <= -11'd95; Sp[752] <= -11'd1019;
Cp[753] <= -11'd89; Sp[753] <= -11'd1020;
Cp[754] <= -11'd83; Sp[754] <= -11'd1020;
Cp[755] <= -11'd76; Sp[755] <= -11'd1021;
Cp[756] <= -11'd70; Sp[756] <= -11'd1021;
Cp[757] <= -11'd64; Sp[757] <= -11'd1021;
Cp[758] <= -11'd58; Sp[758] <= -11'd1022;
Cp[759] <= -11'd51; Sp[759] <= -11'd1022;
Cp[760] <= -11'd45; Sp[760] <= -11'd1022;
Cp[761] <= -11'd39; Sp[761] <= -11'd1023;
Cp[762] <= -11'd33; Sp[762] <= -11'd1023;
Cp[763] <= -11'd26; Sp[763] <= -11'd1023;
Cp[764] <= -11'd20; Sp[764] <= -11'd1023;
Cp[765] <= -11'd14; Sp[765] <= -11'd1023;
Cp[766] <= -11'd7; Sp[766] <= -11'd1023;
Cp[767] <= -11'd1; Sp[767] <= -11'd1023;
Cp[768] <= 11'd4; Sp[768] <= -11'd1023;
Cp[769] <= 11'd11; Sp[769] <= -11'd1023;
Cp[770] <= 11'd17; Sp[770] <= -11'd1023;
Cp[771] <= 11'd23; Sp[771] <= -11'd1023;
Cp[772] <= 11'd29; Sp[772] <= -11'd1023;
Cp[773] <= 11'd36; Sp[773] <= -11'd1023;
Cp[774] <= 11'd42; Sp[774] <= -11'd1023;
Cp[775] <= 11'd48; Sp[775] <= -11'd1022;
Cp[776] <= 11'd55; Sp[776] <= -11'd1022;
Cp[777] <= 11'd61; Sp[777] <= -11'd1022;
Cp[778] <= 11'd67; Sp[778] <= -11'd1021;
Cp[779] <= 11'd73; Sp[779] <= -11'd1021;
Cp[780] <= 11'd80; Sp[780] <= -11'd1020;
Cp[781] <= 11'd86; Sp[781] <= -11'd1020;
Cp[782] <= 11'd92; Sp[782] <= -11'd1019;
Cp[783] <= 11'd98; Sp[783] <= -11'd1019;
Cp[784] <= 11'd105; Sp[784] <= -11'd1018;
Cp[785] <= 11'd111; Sp[785] <= -11'd1017;
Cp[786] <= 11'd117; Sp[786] <= -11'd1017;
Cp[787] <= 11'd123; Sp[787] <= -11'd1016;
Cp[788] <= 11'd130; Sp[788] <= -11'd1015;
Cp[789] <= 11'd136; Sp[789] <= -11'd1014;
Cp[790] <= 11'd142; Sp[790] <= -11'd1014;
Cp[791] <= 11'd148; Sp[791] <= -11'd1013;
Cp[792] <= 11'd155; Sp[792] <= -11'd1012;
Cp[793] <= 11'd161; Sp[793] <= -11'd1011;
Cp[794] <= 11'd167; Sp[794] <= -11'd1010;
Cp[795] <= 11'd173; Sp[795] <= -11'd1009;
Cp[796] <= 11'd179; Sp[796] <= -11'd1008;
Cp[797] <= 11'd186; Sp[797] <= -11'd1006;
Cp[798] <= 11'd192; Sp[798] <= -11'd1005;
Cp[799] <= 11'd198; Sp[799] <= -11'd1004;
Cp[800] <= 11'd204; Sp[800] <= -11'd1003;
Cp[801] <= 11'd210; Sp[801] <= -11'd1002;
Cp[802] <= 11'd216; Sp[802] <= -11'd1000;
Cp[803] <= 11'd223; Sp[803] <= -11'd999;
Cp[804] <= 11'd229; Sp[804] <= -11'd998;
Cp[805] <= 11'd235; Sp[805] <= -11'd996;
Cp[806] <= 11'd241; Sp[806] <= -11'd995;
Cp[807] <= 11'd247; Sp[807] <= -11'd993;
Cp[808] <= 11'd253; Sp[808] <= -11'd992;
Cp[809] <= 11'd259; Sp[809] <= -11'd990;
Cp[810] <= 11'd265; Sp[810] <= -11'd988;
Cp[811] <= 11'd271; Sp[811] <= -11'd987;
Cp[812] <= 11'd277; Sp[812] <= -11'd985;
Cp[813] <= 11'd283; Sp[813] <= -11'd983;
Cp[814] <= 11'd290; Sp[814] <= -11'd982;
Cp[815] <= 11'd296; Sp[815] <= -11'd980;
Cp[816] <= 11'd302; Sp[816] <= -11'd978;
Cp[817] <= 11'd308; Sp[817] <= -11'd976;
Cp[818] <= 11'd314; Sp[818] <= -11'd974;
Cp[819] <= 11'd320; Sp[819] <= -11'd972;
Cp[820] <= 11'd325; Sp[820] <= -11'd970;
Cp[821] <= 11'd331; Sp[821] <= -11'd968;
Cp[822] <= 11'd337; Sp[822] <= -11'd966;
Cp[823] <= 11'd343; Sp[823] <= -11'd964;
Cp[824] <= 11'd349; Sp[824] <= -11'd962;
Cp[825] <= 11'd355; Sp[825] <= -11'd960;
Cp[826] <= 11'd361; Sp[826] <= -11'd958;
Cp[827] <= 11'd367; Sp[827] <= -11'd955;
Cp[828] <= 11'd373; Sp[828] <= -11'd953;
Cp[829] <= 11'd379; Sp[829] <= -11'd951;
Cp[830] <= 11'd384; Sp[830] <= -11'd948;
Cp[831] <= 11'd390; Sp[831] <= -11'd946;
Cp[832] <= 11'd396; Sp[832] <= -11'd944;
Cp[833] <= 11'd402; Sp[833] <= -11'd941;
Cp[834] <= 11'd408; Sp[834] <= -11'd939;
Cp[835] <= 11'd413; Sp[835] <= -11'd936;
Cp[836] <= 11'd419; Sp[836] <= -11'd934;
Cp[837] <= 11'd425; Sp[837] <= -11'd931;
Cp[838] <= 11'd431; Sp[838] <= -11'd928;
Cp[839] <= 11'd436; Sp[839] <= -11'd926;
Cp[840] <= 11'd442; Sp[840] <= -11'd923;
Cp[841] <= 11'd448; Sp[841] <= -11'd920;
Cp[842] <= 11'd453; Sp[842] <= -11'd917;
Cp[843] <= 11'd459; Sp[843] <= -11'd915;
Cp[844] <= 11'd465; Sp[844] <= -11'd912;
Cp[845] <= 11'd470; Sp[845] <= -11'd909;
Cp[846] <= 11'd476; Sp[846] <= -11'd906;
Cp[847] <= 11'd481; Sp[847] <= -11'd903;
Cp[848] <= 11'd487; Sp[848] <= -11'd900;
Cp[849] <= 11'd492; Sp[849] <= -11'd897;
Cp[850] <= 11'd498; Sp[850] <= -11'd894;
Cp[851] <= 11'd503; Sp[851] <= -11'd891;
Cp[852] <= 11'd509; Sp[852] <= -11'd888;
Cp[853] <= 11'd514; Sp[853] <= -11'd885;
Cp[854] <= 11'd520; Sp[854] <= -11'd882;
Cp[855] <= 11'd525; Sp[855] <= -11'd878;
Cp[856] <= 11'd530; Sp[856] <= -11'd875;
Cp[857] <= 11'd536; Sp[857] <= -11'd872;
Cp[858] <= 11'd541; Sp[858] <= -11'd869;
Cp[859] <= 11'd546; Sp[859] <= -11'd865;
Cp[860] <= 11'd552; Sp[860] <= -11'd862;
Cp[861] <= 11'd557; Sp[861] <= -11'd858;
Cp[862] <= 11'd562; Sp[862] <= -11'd855;
Cp[863] <= 11'd568; Sp[863] <= -11'd851;
Cp[864] <= 11'd573; Sp[864] <= -11'd848;
Cp[865] <= 11'd578; Sp[865] <= -11'd844;
Cp[866] <= 11'd583; Sp[866] <= -11'd841;
Cp[867] <= 11'd588; Sp[867] <= -11'd837;
Cp[868] <= 11'd593; Sp[868] <= -11'd834;
Cp[869] <= 11'd599; Sp[869] <= -11'd830;
Cp[870] <= 11'd604; Sp[870] <= -11'd826;
Cp[871] <= 11'd609; Sp[871] <= -11'd823;
Cp[872] <= 11'd614; Sp[872] <= -11'd819;
Cp[873] <= 11'd619; Sp[873] <= -11'd815;
Cp[874] <= 11'd624; Sp[874] <= -11'd811;
Cp[875] <= 11'd629; Sp[875] <= -11'd807;
Cp[876] <= 11'd634; Sp[876] <= -11'd803;
Cp[877] <= 11'd639; Sp[877] <= -11'd800;
Cp[878] <= 11'd644; Sp[878] <= -11'd796;
Cp[879] <= 11'd648; Sp[879] <= -11'd792;
Cp[880] <= 11'd653; Sp[880] <= -11'd788;
Cp[881] <= 11'd658; Sp[881] <= -11'd784;
Cp[882] <= 11'd663; Sp[882] <= -11'd780;
Cp[883] <= 11'd668; Sp[883] <= -11'd775;
Cp[884] <= 11'd672; Sp[884] <= -11'd771;
Cp[885] <= 11'd677; Sp[885] <= -11'd767;
Cp[886] <= 11'd682; Sp[886] <= -11'd763;
Cp[887] <= 11'd687; Sp[887] <= -11'd759;
Cp[888] <= 11'd691; Sp[888] <= -11'd755;
Cp[889] <= 11'd696; Sp[889] <= -11'd750;
Cp[890] <= 11'd700; Sp[890] <= -11'd746;
Cp[891] <= 11'd705; Sp[891] <= -11'd742;
Cp[892] <= 11'd710; Sp[892] <= -11'd737;
Cp[893] <= 11'd714; Sp[893] <= -11'd733;
Cp[894] <= 11'd719; Sp[894] <= -11'd729;
Cp[895] <= 11'd723; Sp[895] <= -11'd724;
Cp[896] <= 11'd727; Sp[896] <= -11'd720;
Cp[897] <= 11'd732; Sp[897] <= -11'd715;
Cp[898] <= 11'd736; Sp[898] <= -11'd711;
Cp[899] <= 11'd741; Sp[899] <= -11'd706;
Cp[900] <= 11'd745; Sp[900] <= -11'd702;
Cp[901] <= 11'd749; Sp[901] <= -11'd697;
Cp[902] <= 11'd753; Sp[902] <= -11'd692;
Cp[903] <= 11'd758; Sp[903] <= -11'd688;
Cp[904] <= 11'd762; Sp[904] <= -11'd683;
Cp[905] <= 11'd766; Sp[905] <= -11'd678;
Cp[906] <= 11'd770; Sp[906] <= -11'd674;
Cp[907] <= 11'd774; Sp[907] <= -11'd669;
Cp[908] <= 11'd779; Sp[908] <= -11'd664;
Cp[909] <= 11'd783; Sp[909] <= -11'd659;
Cp[910] <= 11'd787; Sp[910] <= -11'd654;
Cp[911] <= 11'd791; Sp[911] <= -11'd650;
Cp[912] <= 11'd795; Sp[912] <= -11'd645;
Cp[913] <= 11'd799; Sp[913] <= -11'd640;
Cp[914] <= 11'd802; Sp[914] <= -11'd635;
Cp[915] <= 11'd806; Sp[915] <= -11'd630;
Cp[916] <= 11'd810; Sp[916] <= -11'd625;
Cp[917] <= 11'd814; Sp[917] <= -11'd620;
Cp[918] <= 11'd818; Sp[918] <= -11'd615;
Cp[919] <= 11'd822; Sp[919] <= -11'd610;
Cp[920] <= 11'd825; Sp[920] <= -11'd605;
Cp[921] <= 11'd829; Sp[921] <= -11'd600;
Cp[922] <= 11'd833; Sp[922] <= -11'd595;
Cp[923] <= 11'd836; Sp[923] <= -11'd590;
Cp[924] <= 11'd840; Sp[924] <= -11'd584;
Cp[925] <= 11'd844; Sp[925] <= -11'd579;
Cp[926] <= 11'd847; Sp[926] <= -11'd574;
Cp[927] <= 11'd851; Sp[927] <= -11'd569;
Cp[928] <= 11'd854; Sp[928] <= -11'd564;
Cp[929] <= 11'd858; Sp[929] <= -11'd558;
Cp[930] <= 11'd861; Sp[930] <= -11'd553;
Cp[931] <= 11'd864; Sp[931] <= -11'd548;
Cp[932] <= 11'd868; Sp[932] <= -11'd542;
Cp[933] <= 11'd871; Sp[933] <= -11'd537;
Cp[934] <= 11'd874; Sp[934] <= -11'd532;
Cp[935] <= 11'd878; Sp[935] <= -11'd526;
Cp[936] <= 11'd881; Sp[936] <= -11'd521;
Cp[937] <= 11'd884; Sp[937] <= -11'd516;
Cp[938] <= 11'd887; Sp[938] <= -11'd510;
Cp[939] <= 11'd890; Sp[939] <= -11'd505;
Cp[940] <= 11'd893; Sp[940] <= -11'd499;
Cp[941] <= 11'd896; Sp[941] <= -11'd494;
Cp[942] <= 11'd899; Sp[942] <= -11'd488;
Cp[943] <= 11'd902; Sp[943] <= -11'd483;
Cp[944] <= 11'd905; Sp[944] <= -11'd477;
Cp[945] <= 11'd908; Sp[945] <= -11'd472;
Cp[946] <= 11'd911; Sp[946] <= -11'd466;
Cp[947] <= 11'd914; Sp[947] <= -11'd460;
Cp[948] <= 11'd917; Sp[948] <= -11'd455;
Cp[949] <= 11'd920; Sp[949] <= -11'd449;
Cp[950] <= 11'd922; Sp[950] <= -11'd443;
Cp[951] <= 11'd925; Sp[951] <= -11'd438;
Cp[952] <= 11'd928; Sp[952] <= -11'd432;
Cp[953] <= 11'd930; Sp[953] <= -11'd426;
Cp[954] <= 11'd933; Sp[954] <= -11'd421;
Cp[955] <= 11'd935; Sp[955] <= -11'd415;
Cp[956] <= 11'd938; Sp[956] <= -11'd409;
Cp[957] <= 11'd941; Sp[957] <= -11'd403;
Cp[958] <= 11'd943; Sp[958] <= -11'd398;
Cp[959] <= 11'd945; Sp[959] <= -11'd392;
Cp[960] <= 11'd948; Sp[960] <= -11'd386;
Cp[961] <= 11'd950; Sp[961] <= -11'd380;
Cp[962] <= 11'd952; Sp[962] <= -11'd374;
Cp[963] <= 11'd955; Sp[963] <= -11'd368;
Cp[964] <= 11'd957; Sp[964] <= -11'd363;
Cp[965] <= 11'd959; Sp[965] <= -11'd357;
Cp[966] <= 11'd961; Sp[966] <= -11'd351;
Cp[967] <= 11'd964; Sp[967] <= -11'd345;
Cp[968] <= 11'd966; Sp[968] <= -11'd339;
Cp[969] <= 11'd968; Sp[969] <= -11'd333;
Cp[970] <= 11'd970; Sp[970] <= -11'd327;
Cp[971] <= 11'd972; Sp[971] <= -11'd321;
Cp[972] <= 11'd974; Sp[972] <= -11'd315;
Cp[973] <= 11'd976; Sp[973] <= -11'd309;
Cp[974] <= 11'd977; Sp[974] <= -11'd303;
Cp[975] <= 11'd979; Sp[975] <= -11'd297;
Cp[976] <= 11'd981; Sp[976] <= -11'd291;
Cp[977] <= 11'd983; Sp[977] <= -11'd285;
Cp[978] <= 11'd985; Sp[978] <= -11'd279;
Cp[979] <= 11'd986; Sp[979] <= -11'd273;
Cp[980] <= 11'd988; Sp[980] <= -11'd267;
Cp[981] <= 11'd990; Sp[981] <= -11'd261;
Cp[982] <= 11'd991; Sp[982] <= -11'd255;
Cp[983] <= 11'd993; Sp[983] <= -11'd249;
Cp[984] <= 11'd994; Sp[984] <= -11'd242;
Cp[985] <= 11'd996; Sp[985] <= -11'd236;
Cp[986] <= 11'd997; Sp[986] <= -11'd230;
Cp[987] <= 11'd999; Sp[987] <= -11'd224;
Cp[988] <= 11'd1000; Sp[988] <= -11'd218;
Cp[989] <= 11'd1001; Sp[989] <= -11'd212;
Cp[990] <= 11'd1003; Sp[990] <= -11'd206;
Cp[991] <= 11'd1004; Sp[991] <= -11'd199;
Cp[992] <= 11'd1005; Sp[992] <= -11'd193;
Cp[993] <= 11'd1006; Sp[993] <= -11'd187;
Cp[994] <= 11'd1007; Sp[994] <= -11'd181;
Cp[995] <= 11'd1008; Sp[995] <= -11'd175;
Cp[996] <= 11'd1009; Sp[996] <= -11'd169;
Cp[997] <= 11'd1010; Sp[997] <= -11'd162;
Cp[998] <= 11'd1011; Sp[998] <= -11'd156;
Cp[999] <= 11'd1012; Sp[999] <= -11'd150;
Cp[1000] <= 11'd1013; Sp[1000] <= -11'd144;
Cp[1001] <= 11'd1014; Sp[1001] <= -11'd137;
Cp[1002] <= 11'd1015; Sp[1002] <= -11'd131;
Cp[1003] <= 11'd1016; Sp[1003] <= -11'd125;
Cp[1004] <= 11'd1017; Sp[1004] <= -11'd119;
Cp[1005] <= 11'd1017; Sp[1005] <= -11'd112;
Cp[1006] <= 11'd1018; Sp[1006] <= -11'd106;
Cp[1007] <= 11'd1019; Sp[1007] <= -11'd100;
Cp[1008] <= 11'd1019; Sp[1008] <= -11'd94;
Cp[1009] <= 11'd1020; Sp[1009] <= -11'd87;
Cp[1010] <= 11'd1020; Sp[1010] <= -11'd81;
Cp[1011] <= 11'd1021; Sp[1011] <= -11'd75;
Cp[1012] <= 11'd1021; Sp[1012] <= -11'd69;
Cp[1013] <= 11'd1022; Sp[1013] <= -11'd62;
Cp[1014] <= 11'd1022; Sp[1014] <= -11'd56;
Cp[1015] <= 11'd1022; Sp[1015] <= -11'd50;
Cp[1016] <= 11'd1023; Sp[1016] <= -11'd44;
Cp[1017] <= 11'd1023; Sp[1017] <= -11'd37;
Cp[1018] <= 11'd1023; Sp[1018] <= -11'd31;
Cp[1019] <= 11'd1023; Sp[1019] <= -11'd25;
Cp[1020] <= 11'd1023; Sp[1020] <= -11'd18;
Cp[1021] <= 11'd1023; Sp[1021] <= -11'd12;
Cp[1022] <= 11'd1023; Sp[1022] <= -11'd6;
Cp[1023] <= 11'd1024; Sp[1023] <= -11'd0;

end

// Running sums for B* ( c*x, s*x, c*y, s*y )
reg signed [25:0] Cpx;
reg signed [25:0] Spx;
reg signed [25:0] Cpy;
reg signed [25:0] Spy;

// Actual x' and y'
wire [25:0] xp_divd = (Cpx - Spy) >>> 10;
wire [25:0] yp_divd = (Spx + Cpy) >>> 10;

// Index into the 
reg [9:0] theta_i = 0;

// Advance x,y based on pixel clock, update rotation sums,
// update frame counter, and update theta index each frame
always @(posedge clk25)
begin
  if (pix_x < hpixels - 1) begin
    pix_x <= pix_x + 1;
    Cpx <= Cpx + Cp[theta_i];
    Spx <= Spx + Sp[theta_i];
  end
  else
  begin
    // Next line
    pix_x <= 0;
    Cpx <= 0;
    Spx <= 0;

    if (pix_y < vlines - 1) begin
      pix_y <= pix_y + 1;
      Cpy <= Cpy + Cp[theta_i];
      Spy <= Spy + Sp[theta_i];
    end

    else begin
      pix_y <= 0;
      Cpy <= 0;
      Spy <= 0;
      frame_counter <= frame_counter + 1;
      if (frame_counter[0])
        theta_i <= theta_i + 1;
      else
        theta_i <= theta_i;
    end
  end

  // Shift tile data (x,y) indexing by looking up line_shifts data
  // The divide by 4 is just to enlarge tiles which looks nice.
  //
  // (x,y) are not used, but rather (x',y') so rotation also occurs
  shift_x_index = yp_divd[5:0] + frame_counter[5:0];
  shift_x = (xp_divd[5:0] + 16 - line_shifts[ shift_x_index ]) / 4;
  shift_y_index = xp_divd[5:0] + frame_counter[5:0];
  shift_y = (yp_divd[5:0] + 16 - line_shifts[ shift_y_index ]) / 4;
  pix_reg = tile_data[ shift_y[2:0] ][ shift_x[2:0] ];
end

// In this video mode, hsync and vsync are active low when the pulse
// is supposed to take place
assign hsync = (pix_x >= (res_x+hfp) && pix_x < (res_x+hfp+hpulse)) ? 0 : 1;
assign vsync = (pix_y >= (res_y+vfp) && pix_y < (res_y+vfp+vpulse)) ? 0 : 1;

wire pix_on = pix_reg;

always @*
begin
  // first check if we're within vertical active video range
  if (pix_y < res_y && pix_x < res_x)
  begin
    // Some color variation in a kind of checkerboard pattern
    r0 <= (shift_y[3] ^ shift_x[3]) ? pix_on : 0;
    g0 <= ~(shift_y[3] ^ shift_x[3]) ? pix_on : 0;
    b0 <= (shift_y[4] ^ shift_x[4]) ? pix_on : 0;
  end
  else
  begin
    // If we're outside the visible frame, it's important to
    // actually set 0. (My monitor doesn't show anything otherwise)
    r0 <= 0;
    g0 <= 0;
    b0 <= 0;
  end
end

endmodule

